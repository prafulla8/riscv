module \$_DLATCH_N_ (E, D, Q);
//  wire [1023:0] _TECHMAP_DO_ = "simplemap; opt";
  input E, D;
  output Q;
  sky130_fd_sc_hd__dlxtp_1 _TECHMAP_REPLACE_ (
    .D(D),
    .GATE(E),
    .Q(Q)
  );
endmodule

module \$_DLATCH_P_ (E, D, Q);
//  wire [1023:0] _TECHMAP_DO_ = "simplemap; opt";
  input E, D;
  output Q;
  sky130_fd_sc_hd__dlxtp_1 _TECHMAP_REPLACE_ (
    .D(D),
    .GATE(E),
    .Q(Q)
  );
endmodule
